`timescale 1ns/1ns

module test_FSM();
wire [1:0]state;
reg inp;
wire out;
aaaaaa F1(state,inp,out);
initial begin
inp=0;
#5 inp=1;
end

initial begin
#5 inp=0;
#5 inp=1;
#5 inp=0;
#5 inp=1;
end
endmodule
