module practice(a,b,cin,s,cout);

input [3:0] a,b;
input cin;
wire [3:0] w;
output [3:0] s;
output cout;

full_adder f1(a[0],b[0],cin,s[0],w[0]);
full_adder f2(a[1],b[1],w[0],s[1],w[1]);
full_adder f3(a[2],b[2],w[1],s[2],w[2]);
full_adder f4(a[3],b[3],w[2],s[3],w[3]);

assign cout = w[3];

endmodule
