




`timescale 1ns/1ns

module test_seven_segment();
	reg [2:0]a;
	wire [15:0]out;
	seven_segment F1(a,out);
	
	initial begin 
	a = 3'b001;
	#20 a = 3'b010;
	#20 a = 3'b011;
	#20 a = 3'b100;
	#10 $finish;
	end
	
	
 	
endmodule 