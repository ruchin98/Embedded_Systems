module not_gate (a,b);

	input a;
	output b;
	assign b=~a;
	
endmodule 
